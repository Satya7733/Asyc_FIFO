package AFIFO_Pkg;
  `include "AFIFO_Transaction.sv"
  `include "AFIFO_Generator.sv"
  `include "AFIFO_Driver.sv"
  `include "AFIFO_Monitor.sv"
  `include "AFIFO_Scoreboard.sv"
  `include "AFIFO_Environment.sv"
endpackage
