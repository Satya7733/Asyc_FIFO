class driver;


endclass
