`include "wr_intf.sv"
`include "rd_intf.sv"
`include "trans.sv"

