//  `include "FIFO.sv"
//  `include "uvm_AFIFO_sequence_item.sv"
//  `include "uvm_AFIFO_sequence.sv"
//  `include "uvm_AFIFO_driver.sv"
//  `include "uvm_AFIFO_monitor.sv"
//  `include "uvm_AFIFO_scoreboard.sv"
//
