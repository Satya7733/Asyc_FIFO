//imports
import AFIFO_Pkg::*;

//class
class AFIFO_Monitor #(parameter DSIZE = 8);

//Transaction class initialize
AFIFO_Transaction tr_mon2scb;

// Handle
virtual AFIFO_Interface vif_mon;

//Mailbox mon to sco
mailbox #(AFIFO_Transaction) mbx_mon2sco;

//Constructor
function new(mailbox #(AFIFO_Transaction) mbx_mon2sco);
 this.mbx_mon2sco = mbx_mon2sco;
endfunction

//Event
event mon_done;
//Task
task run();
 tr_mon2scb = new();
forever begin
 /*   
 @(posedge vif.rd_clk); 
 if(vif.rd_inc && !vif.rd_empty) begin
 mbx_mon2sco.put(vif.rd_data);
  $display("[MON]:----------------------------------------");
 $display("[MON]: MBX DATA SENT TO SCO %0d ", vif.rd_data);
 
 end
   $display("[MON]:----------------------------------------");
 if(vif.rd_empty) $display("[MON] : READ EMPTY, Nothing to read in FIFO Mem ");
 if(vif.wr_full) $display("[MON] : WRITE FULL, Full FIFO Mem ");
  $display("[MON]:----------------------------------------");
 */

 @(posedge vif_mon.rd_inc or posedge vif_mon.wr_inc); 
if(vif_mon.rd_inc || vif_mon.rd_empty || vif_mon.wr_full || ~vif_mon.rd_rst || ~vif_mon.rd_rst || vif_mon.wr_inc) begin 
$display("[MON]:Entered Loop sending Tr class");
//5ns
 tr_mon2scb.rd_data <= vif_mon.rd_data;
 tr_mon2scb.wr_inc <= vif_mon.wr_inc;
 tr_mon2scb.rd_inc <= vif_mon.rd_inc;
 tr_mon2scb.wr_rst <= vif_mon.wr_rst;
 tr_mon2scb.rd_rst <= vif_mon.rd_rst;
 tr_mon2scb.rd_empty <= vif_mon.rd_empty;
 tr_mon2scb.wr_full <= vif_mon.wr_full;
$display("[MON]: rd_inc = %d, wr_inc = %d", tr_mon2scb.rd_inc, tr_mon2scb.wr_inc);
if(vif_mon.rd_inc)$display("[MON]: MBX DATA SENT TO SCO %0d ", tr_mon2scb.rd_data);
 mbx_mon2sco.put(tr_mon2scb);
 if(vif_mon.rd_inc)$display("[MON]: MBX DATA SENT TO SCO %0d ", tr_mon2scb.rd_data);
 ->mon_done;
if(vif_mon.rd_inc)$display("[MON]: MBX DATA SENT TO SCO %0d ", tr_mon2scb.rd_data);
//$display("[MON]:----------------------------------------");
end
end

endtask

endclass
