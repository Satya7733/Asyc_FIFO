class transaction;

rand bit [DATASIZE-1:0] idata;
rand bit 		wren;
rand bit 		rden;
bit 			wrst;
bit			rrst;

endclass : transaction

