interface AFIFO_Interface #(parameter DSIZE = 8,parameter ASIZE = 4);
	logic [DSIZE-1:0] rd_data;
	logic [DSIZE-1:0] wr_data;
	logic wr_full;
	logic rd_empty;
	logic wr_inc;
	logic rd_inc;
	logic wr_clk;
	logic rd_clk;
	logic wr_rst;
	logic rd_rst;
endinterface
