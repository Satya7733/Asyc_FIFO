
`include "uvm_macros.svh"
import uvm_pkg::*;
import uvm_AFIFO_agent_pkg::*;

typedef uvm_sequencer#(uvm_AFIFO_Wr_sequence_item) write_sequencer;

