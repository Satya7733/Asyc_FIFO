
`include "uvm_macros.svh"
import uvm_pkg::*;

//`include "uvm_AFIFO_agent_pkg.sv"
import uvm_AFIFO_agent_pkg::*;



typedef uvm_sequencer#(uvm_AFIFO_Rd_sequence_item) read_sequencer;

